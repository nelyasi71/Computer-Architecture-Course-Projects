`define BEQ 3'b000
`define BNE 3'b001
`define BLT 3'b010
`define BGE 3'b011

module BranchController(input [2:0] func3, input branch, zero, neg, output reg w);
    
    always @(func3, zero, neg, branch) begin
        case(func3)
            `BEQ   : w <= branch & zero;
            `BNE   : w <= branch & ~zero;
            `BLT   : w <= branch & neg;
            `BGE   : w <= branch & (zero | ~neg);
            default: w <= 1'b0;
        endcase
    end

endmodule